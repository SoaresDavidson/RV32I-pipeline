module control(
    
);
endmodule