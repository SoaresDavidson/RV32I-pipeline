module BranchDecider (
  input  wire [6:0] opcode,
  input  wire [2:0] funct3,
  input  wire [31:0] rs1,
  input  wire [31:0] rs2,
  input  wire [11:0] imm,
  output reg  Branch,
  output reg  [11:0] Deviation
);
  always @(*) begin
    // valores padrão
    Branch    = 1'b0;
    Deviation = 12'b0;

    if (opcode == 7'b1100011) begin
      case (funct3)
        3'b000: Branch = (rs1 == rs2);   // BEQ
        3'b001: Branch = (rs1 != rs2);   // BNE
        3'b100: Branch = (rs1 < rs2);    // BLT
        3'b101: Branch = (rs1 >= rs2);   // BGE
        3'b110: Branch = ($signed(rs1) < $signed(rs2)) // BLT signed
        3'b111: Branch = ($signed(rs1) >= $signed(rs2)) // BGE signed
        default: Branch = 1'b0;
      endcase

      if (Branch)
        Deviation = imm;
    end
  end
endmodule