module R232i;
  
  reg [31:0]A;
  reg [31:0]B;
  wire [31:0]C;
  wire z;
  reg [1:0]sel;

  ULA dut ( .A (A),
            .B (B),
				.C (C),
				.z (z),
				.sel (sel)
	);
	
endmodule